// Background image display

module background
	(
		CLOCK_50,						//	On Board 50 MHz
		KEY,							//	Push Button[0:0]
		VGA_CLK,   						//	VGA Clock
		VGA_HS,							//	VGA H_SYNC
		VGA_VS,							//	VGA V_SYNC
		VGA_BLANK,						//	VGA BLANK
		VGA_SYNC,						//	VGA SYNC
		VGA_R,   						//	VGA Red[9:0]
		VGA_G,	 						//	VGA Green[9:0]
		VGA_B	  						//	VGA Blue[9:0]
	);

	input	CLOCK_50;				//	50 MHz
	input	[0:0] KEY;				//	Button[0:0]
	output	VGA_CLK;   				//	VGA Clock
	output	VGA_HS;					//	VGA H_SYNC
	output	VGA_VS;					//	VGA V_SYNC
	output	VGA_BLANK;				//	VGA BLANK
	output	VGA_SYNC;				//	VGA SYNC
	output	[9:0] VGA_R;   			//	VGA Red[9:0]
	output	[9:0] VGA_G;	 		//	VGA Green[9:0]
	output	[9:0] VGA_B;   			//	VGA Blue[9:0]
	
	wire resetn, gnd;
	reg [0:0] reg_gnd;
	assign resetn = KEY[0];
	assign gnd = reg_gnd;
	
	// Create the color, x, y and writeEn wires that are inputs to the controller.

	wire [2:0] color;
	reg [7:0] x;
	reg [6:0] y;
	assign color = 3'd0;
	
	always@(posedge CLOCK_50 or negedge resetn)begin
		if (!resetn)begin
			x <= 8'd0;
			y <= 7'd0;
			reg_gnd <= 1'b0;
		end
		else begin
			if ((x == 8'd2) && (y == 7'd2))
				reg_gnd <= 1'b0;
			else begin
				x <= (x == 8'd2)? (8'd0) : (x + 8'd1);
				y <= (x == 8'd2)? (y + 7'd1) : y;
				reg_gnd <= 1'b1;
			end
		end
	end
	
	// Create an Instance of a VGA controller - "There can be only one!"
	// Define the number of colours as well as the initial background
	// image file (.MIF) for the controller.
	vga_adapter VGA(
			.resetn(resetn),
			.clock(CLOCK_50),
			.colour(color),
			.x(x),
			.y(y),
			.plot(gnd),
			/* Signals for the DAC to drive the monitor. */
			.VGA_R(VGA_R),
			.VGA_G(VGA_G),
			.VGA_B(VGA_B),
			.VGA_HS(VGA_HS),
			.VGA_VS(VGA_VS),
			.VGA_BLANK(VGA_BLANK),
			.VGA_SYNC(VGA_SYNC),
			.VGA_CLK(VGA_CLK));
		defparam VGA.RESOLUTION = "160x120";
		defparam VGA.MONOCHROME = "FALSE";
		defparam VGA.BITS_PER_COLOUR_CHANNEL = 1;
		defparam VGA.BACKGROUND_IMAGE = "display.mif";
		
endmodule
